`timescale 1ns / 1ps

/*
 * Testbench for pdpm memory part, i.e. the block diagram
 */

module pdpm_mem_tb(

    );
endmodule
