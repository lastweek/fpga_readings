module hello_world;

initial begin
	$display("Hello world to where?");
	$display("And this is hacked by simulator?");
end

endmodule
